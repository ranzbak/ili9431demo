/**
 * PLL configuration
 *
 * This Verilog module was generated automatically
 * using the icepll tool from the IceStorm project.
 * Use at your own risk.
 *
 * Given input frequency:        16.000 MHz
 * Requested output frequency:   21.477 MHz
 * Achieved output frequency:    21.500 MHz
 */

module pll(
    input  clock_in,
    output clock_out,
    output locked
);

    // 12 MHz in
    // 16 MHz out

    SB_PLL40_CORE #(
    .FEEDBACK_PATH("SIMPLE"),
    .DIVR(4'b0000), // DIVR =  0
    .DIVF(7'b1010100), // DIVF = 42
    .DIVQ(3'b101), // DIVQ =  5
    .FILTER_RANGE(3'b001) // FILTER_RANGE = 1
    ) uut (
        .LOCK(locked),
        .RESETB(1'b1),
        .BYPASS(1'b0),
        .REFERENCECLK(clock_in),
        .PLLOUTCORE(clock_out)
    );

endmodule